# This is the Swedish language file for ImageViewer.

# The structure of the file is as follows:

# A line starting with "#" is interpreted as a comment.

# A valid non comment line may look like "file = Arkiv" where "file" is the variable, = the
# separator and "Arkiv" is the value of the variable, in this case the Swedish word for file.

# There might be whitespaces or tabs in between the variable and the "=". Any whitespace
# or other character after the value of the variable will be trimmed away.

# For more information regarding the rules for the syntax of this file please visit:
# http://java.sun.com/javase/6/docs/api/java/util/Properties.html

# This file was created: by Fredrik M�ller 2009-08-20
# This file was updated: 

##############################################################################################################
# I M A G E  V I E W E R                                                                                     #
##############################################################################################################
imageviewer.button.back.toolTip                         = F�reg�ende (V�nsterpil) 
imageviewer.button.forward.toolTip                      = N�sta (H�gerpil) 
imageviewer.button.automaticAdjustToWindowSize.toolTip  = Automatisk anpassning till f�nsterstorlek (Alt + C) 
imageviewer.button.automaticAdjustToWindowSize.mnemonic = C
imageviewer.button.adjustToWindowSize.toolTip           = Anpassa till f�nsterstorlek (Alt + A) 
imageviewer.button.adjustToWindowSize.mnemonic          = A
imageviewer.button.help.toolTip                         = Hj�lp (Alt + H) 
imageviewer.button.help.mnemonic                        = H
imageviewer.button.rotateLeft.toolTip                   = Rotera bild v�nster (Alt + V�nsterpil)
imageviewer.button.rotateRight.toolTip                  = Rotera bild h�ger (Alt + H�gerpil)
imageviewer.button.rotateAutomatic                      = Rotera bild automatiskt (Alt + Pil Upp)

imageviewer.popupmenu.back.text               = (Alt-Z) F�reg�ende
imageviewer.popupmenu.forward.text            = (Alt-X) N�sta
imageviewer.popupmenu.adjustToWindowSize.text = (Alt-A) Anpassa till f�nsterstorlek

imageviewer.statusbar.pathToPicture    = S�kv�g till bildfilen
imageviewer.statusbar.sizeLabel        = S:
imageviewer.statusbar.sizeLabelImage   = Bildstorlek i 
imageviewer.statusbar.widthLabel       = B:
imageviewer.statusbar.widthLabelImage  = Bildbredd i pixlar
imageviewer.statusbar.heightLabel      = H:
imageviewer.statusbar.heightLabelImage = Bildh�jd i pixlar

##############################################################################################################
# M E T A  D A T A  P A N E L                                                                                #
##############################################################################################################
metadatapanel.titleDefaultText     = METADATA F�R BILD:
metadatapanel.tableheader.type     = TYP
metadatapanel.tableheader.property = EGENSKAP
metadatapanel.tableheader.value    = V�RDE

##############################################################################################################
# I M A G E  S E A R C H  R E S U L T  V I E W E R                                                                                     #
##############################################################################################################
imagesearchresultviewer.title = S�kresultat
imagesearchresultviewer.menuitem.selectAll = Markera alla bilder
imagesearchresultviewer.menuitem.deSelectAll = Avmarkera alla markerade bilder
imagesearchresultviewer.menuitem.addSelectedImagesToViewList = L�gg valda bilder till bildlistan
imagesearchresultviewer.menuitem.copySelectedImagesToSystemClipboard = Kopiera valda bilder till systemets urklippshanterare
imagesearchresultviewer.menuitem.copyAllImagesToSystemClipboard = Kopiera alla bilder till systemets urklippshanterare
imagesearchresultviewer.statusMessage.amountOfImagesInSearchResult = Antal bilder i s�kresultatet