# This is the Swedish language file for the image statistics viewer strings.

# The structure of the file is as follows:

# A line starting with "#" is interpreted as a comment.

# A valid non comment line may look like "file = Arkiv" where "file" is the variable, = the
# separator and "Arkiv" is the value of the variable, in this case the Swedish word for file.

# There might be whitespaces or tabs in between the variable and the "=". Any whitespace
# or other character after the value of the variable will be trimmed away.

# For more information regarding the rules for the syntax of this file please visit:
# http://java.sun.com/javase/6/docs/api/java/util/Properties.html

##############################################################################################################
# C O M M O N  T E X T S                                                                                     #
##############################################################################################################
imagestatisticsviewer.chart.title.prefix = Antal bilder per: 
imagestatisticsviewer.chart.valueAxisLabel = antal bilder

##############################################################################################################
# T A B  S P E C I F I C  T E X T                                                                            #
##############################################################################################################
imagestatisticsviewer.chart.weekday.title = Veckodag
imagestatisticsviewer.chart.fnumber.title = Bländartal
imagestatisticsviewer.chart.exposuretime.title = Exponeringstid
imagestatisticsviewer.chart.iso.title = ISO
imagestatisticsviewer.chart.imagesize.title = Bildstorlek
imagestatisticsviewer.chart.second.title = Sekund
imagestatisticsviewer.chart.minute.title = Minut
imagestatisticsviewer.chart.hour.title = Timme
imagestatisticsviewer.chart.dayinmonth.title = Dag i månad
imagestatisticsviewer.chart.year.title = År
imagestatisticsviewer.chart.cameramodel.title = Kameramodell