category.categoriesModel.create.error = Kan inte ladda kategorier.\nJavaPEG kommer att avslutas\n\nSe loggfil för detaljer.
category.categoriesModel.store.error  = Kan inte spara kategorier.\nJavaPEG kommer att avslutas\n\nSe loggfil för detaljer.

category.categoriesModel.repositoryExists       = Bilddatabassökväg existerar.
category.categoriesModel.repositoryNotExists    = Bilddatabassökväg existerar inte.
category.categoriesModel.repositoryNotAvailable = Bilddatabassökväg inte tillgänglig.

category.metadatavalue.selection.mode   = URVALSMETOD
category.metadatavalue.selection.values = VÄRDEN

category.enterNameForNewCategory    = Ange ett namn för den nya kategorin
category.enterNameForNewSubCategory = Ange ett namn för den nya underkategorin
category.enterNewNameForCategory    = Ange ett nytt namn för den kategorin:
categrory.rename                    = Byt namn på kategori

category.errormessage.categoryNameCanNotStartWithSpace = Kategorinamnet kan inte börja med ett mellanslag:
category.errormessage.categoryNameAlreadyExistsInScope = existerar redan som en kategori i vald kontext, välj ett annat namn

category.addToImageRepositoryHeader = Lägg till bild(er) till bilddatabas?
category.addToImageRepositoryQuestionPartOne = Lägg till bild(erna) i katalog:
category.addToImageRepositoryQuestionPartTwo = till bilddatabasen?

category.rememberMySelection = Kom ihåg mitt val (Kan ändras i Inställningarna)

category.mineCategoriesTab = Mina