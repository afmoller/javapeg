# This is the Swedish language file for the Image Merge Functionality.

# The structure of the file is as follows:

# A line starting with "#" is interpreted as a comment.

# A valid non comment line may look like "file = Arkiv" where "file" is the variable, = the
# separator and "Arkiv" is the value of the variable, in this case the Swedish word for file.

# There might be whitespaces or tabs in between the variable and the "=". Any whitespace
# or other character after the value of the variable will be trimmed away.

# For more information regarding the rules for the syntax of this file please visit:
# http://java.sun.com/javase/6/docs/api/java/util/Properties.html

imagemerge.gui.title = KATALOGER ATT SLÅ SAMMAN
imagemerge.gui.conflict.viewer.title = Sammanslagningskonfliktsvisare

imagemerge.processlog.title = PROCESSLOGG

imagemerge.tooltip.directories.remove   = Ta bort vald katalog
imagemerge.tooltip.directories.add      = Lägg till visad katalog
imagemerge.tooltip.process.merge.start  = Slå samman bilder från de valda katalogerna
imagemerge.tooltip.process.merge.cancel = Avbryt sammanslagningsprocessen

imagemerge.process.md5Sum.calculated = MD5 summa beräknad (%s) för fil: %s (%s millisekunder)

imagemerge.process.started        = Sammanslagningsprocess startad
imagemerge.process.aborted        = Sammanslagningsprocess avbruten
imagemerge.process.done           = Sammanslagningsprocessen tog: %s sekunder
imagemerge.process.done.cancelled = Sammanslagningsprocessen avbröts efter: %s sekunder
imagemerge.process.done.popup           = Sammanslagning färdig
imagemerge.process.done.popup.cancelled = Sammanslagning avbruten


imagemerge.process.destinationdirectory.created     = Destinationskatalog skapad:
imagemerge.process.destinationdirectory.not.created = Destinationskatalog kunde inte skapas:

imagemerge.process.images.searching       = Letar efter JPEG-filer i valda kataloger
imagemerge.process.images.searching.found = JPEG-filer funna i katalog:

imagemerge.process.images.copy.started  = Kopieringsprocessen startad
imagemerge.process.images.copy.image    = Fil: %s kopierades till destinationskatalogen med namnet:
imagemerge.process.images.copy.finished = Kopieringsprocessen avslutad

imagemerge.conflict.viewer = Bild: %s valdes i bildkonfliktsvisaren
