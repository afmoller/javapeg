###################################################################################################
# This is the Swedish language file for HelpViewer.
#
# The structure of the file is as follows:
#
# A line starting with "#" is interpreted as a comment.
#
# A valid non comment line may look like "file = Arkiv" where "file" is the variable, = the
# separator and "Arkiv" is the value of the variable, in this case the Swedish word for file.
#
# There might be whitespaces or tabs in between the variable and the "=". Any whitespace
# or other character after the value of the variable will be trimmed away.
#
# For more information regarding the rules for the syntax of this file please visit:
# http://java.sun.com/javase/6/docs/api/java/util/Properties.html
###################################################################################################
helpViewerGUI.window.locationError = Kunde inte sätta fönsterposition enligt konfigurationen. Se loggfil för detaljer.
helpViewerGUI.window.title         = Hjälp
helpViewerGUI.errorMessage         = Kunde inte ladda hjälpfil, se loggfil för detaljer.

helpViewerGUI.tree.content                    = Innehåll
helpViewerGUI.tree.programHelpOverView        = PROGRAMBESKRIVNING
helpViewerGUI.tree.programHelpMerge           = SLÅ IHOP BILDER
helpViewerGUI.tree.programHelpRename          = BYT NAMN PÅ BILDER
helpViewerGUI.tree.programHelpViewImages      = VISA BILDER
helpViewerGUI.tree.programHelpImagesTag       = TAGGA BILDER
helpViewerGUI.tree.programHelpImagesSearch    = SÖK BILDER
helpViewerGUI.tree.programHelpImageViewer     = BILDVISARE
helpViewerGUI.tree.programHelpImageResizer    = BILDSTORLEKSÄNDRARE
helpViewerGUI.tree.programHelpOverviewCreator = SKAPA TUMNAGELÖVERSIKT
helpViewerGUI.tree.versionInformation         = VERSIONSINFORMATION
helpViewerGUI.tree.references                 = REFERENSER / TACK TILL
helpViewerGUI.tree.configuration              = Inställningar
helpViewerGUI.tree.logging                    = LOGGNING
helpViewerGUI.tree.updates                    = UPPDATERINGAR
helpViewerGUI.tree.rename                     = NAMNBYTE
helpViewerGUI.tree.language                   = SPRÅK
helpViewerGUI.tree.thumbnail                  = TUMNAGEL
helpViewerGUI.tree.tag                        = TAGGAR
helpViewerGUI.tree.functionality              = Funktionalitet
helpViewerGUI.tree.problems                   = Problem
helpViewerGUI.tree.corrupt                    = BILDDATABAS KORRUPT
helpViewerGUI.tree.inconsistent               = BILDDATABAS INKONSISTENT