# This is the Swedish language file for the Image repository part of JavaPEG.

# The structure of the file is as follows:

# A line starting with "#" is interpreted as a comment.

# A valid non comment line may look like "file = Arkiv" where "file" is the variable, = the
# separator and "Arkiv" is the value of the variable, in this case the Swedish word for file.

# There might be whitespaces or tabs in between the variable and the "=". Any whitespace
# or other character after the value of the variable will be trimmed away.

# For more information regarding the rules for the syntax of this file please visit:
# http://java.sun.com/javase/6/docs/api/java/util/Properties.html

imagerepository.addDirectoryToAllwaysAddAutomaticallyList.label = L�gg till katalog till listan av kataloger d�r bilder l�ggs till i bilddatabasen automatiskt
imagerepository.addDirectoryToNeverAddAutomaticallyList.label   = L�gg till katalog till listan av kataloger d�r bilder inte skall l�ggas till automatiskt till bilddatabasen

imagerepository.repositoryfile.corrupt.1 = The repository file is corrupt
imagerepository.repositoryfile.corrupt.2 = The corrupt repository file was succesfully backed up to the file:
imagerepository.repositoryfile.corrupt.3 = Could not back up the repository file. Content is written to JavaPEG log file
imagerepository.repositoryfile.corrupt.4 = Repository file restored to default
imagerepository.repositoryfile.corrupt.5 = Could not restore the repository file to default
imagerepository.repositoryfile.corrupt.6 = Please add the following content manually to the repository file:
imagerepository.repositoryfile.corrupt.7 = Content start:
imagerepository.repositoryfile.corrupt.8 = Could not fetch content
imagerepository.repositoryfile.corrupt.9 = Content end:
imagerepository.repositoryfile.corrupt.10 = See JavaPEG log file for details

imagerepository.model.store.error  = Could not save image repository, see log file for details
imagerepository.model.create.error = Could not load image repository, see log file for details

imagerepository.directory.added                = Selected directory is part of the image repository database
imagerepository.directory.added.writeprotected = Selected directory is part of the image repository database, but the database file is write protected
imagerepository.directory.not.added            = Selected directory is not part of the image repository database