# This is the Swedish language file for the Image repository part of JavaPEG.

# The structure of the file is as follows:

# A line starting with "#" is interpreted as a comment.

# A valid non comment line may look like "file = Arkiv" where "file" is the variable, = the
# separator and "Arkiv" is the value of the variable, in this case the Swedish word for file.

# There might be whitespaces or tabs in between the variable and the "=". Any whitespace
# or other character after the value of the variable will be trimmed away.

# For more information regarding the rules for the syntax of this file please visit:
# http://java.sun.com/javase/6/docs/api/java/util/Properties.html

imagerepository.addDirectoryToAllwaysAddAutomaticallyList.label = L�gg till katalog till listan av kataloger d�r bilder l�ggs till i bilddatabasen automatiskt
imagerepository.addDirectoryToNeverAddAutomaticallyList.label   = L�gg till katalog till listan av kataloger d�r bilder inte skall l�ggas till automatiskt till bilddatabasen

imagerepository.repositoryfile.corrupt.1 = Bilddatabasfilen �r korrupt
imagerepository.repositoryfile.corrupt.2 = Den korrupta bilddatabasfilen s�kerhetskopierades korrekt:
imagerepository.repositoryfile.corrupt.3 = Kunde inte s�kerhetskopiera bilddatabasfilen. Inneh�llet har skrivits till JavaPEGs loggfil
imagerepository.repositoryfile.corrupt.4 = Bilddatabasfilen har �terst�llts till ursprungligt skick.
imagerepository.repositoryfile.corrupt.5 = Kunde inte �terst�lla bilddatabasfilen till ursprungligt skick
imagerepository.repositoryfile.corrupt.6 = V�nligen mata inte f�ljande inneh�ll manuellt i bilddatabasen:
imagerepository.repositoryfile.corrupt.7 = Start inneh�ll:
imagerepository.repositoryfile.corrupt.8 = Kunde inte h�mta inneh�ll
imagerepository.repositoryfile.corrupt.9 = Inneh�ll slut:
imagerepository.repositoryfile.corrupt.10 = Se JavaPEGs loggfil f�r detaljer

imagerepository.model.store.error  = Kunde inte spara bilddatabasen, se loggfil f�r detaljer.
imagerepository.model.create.error = Kunde inte �ppna bilddatabasen, se loggfil f�r detaljer.

imagerepository.directory.added                = Vald katalog �r en del av bilddatabasen
imagerepository.directory.added.writeprotected = Vald katalog �r en del av bilddatabasen, men databasfilen �r skrivskyddad
imagerepository.directory.not.added            = Vald katalog �r inte en del av bilddatabasen

imagerepository.directory.already.added.to.allways.add         = har redan blivit tillagd i listan av kataloger f�r vilka\n bilder alltid kommer att l�ggas till automatiskt till bilddatabasen.
imagerepository.directory.already.added.to.never.add           = har redan blivit tillagd i listan av kataloger f�r vilka\n bilder aldrig kommer att l�ggas till automatiskt till bilddatabasen.
imagerepository.directory.is.parent.to.already.added.directory = En underkatalog har redan blivit tillagd i listan av kataloger\n f�r vilka bilder alltid kommer att l�ggas till automatiskt \ntill bilddatabasen eller i listan av kataloger f�r vilka bilder\n aldrig kommer att l�ggas till automatiskt till bilddatabasen.\n\nSe JavaPEGs inst�llningar f�r detaljer.