# This is the Swedish language file for the common strings.

# The structure of the file is as follows:

# A line starting with "#" is interpreted as a comment.

# A valid non comment line may look like "file = Arkiv" where "file" is the variable, = the
# separator and "Arkiv" is the value of the variable, in this case the Swedish word for file.

# There might be whitespaces or tabs in between the variable and the "=". Any whitespace
# or other character after the value of the variable will be trimmed away.

# For more information regarding the rules for the syntax of this file please visit:
# http://java.sun.com/javase/6/docs/api/java/util/Properties.html

common.button.ok.label = Ok
common.button.apply.label = Verkst�ll
common.button.cancel.label = Avbryt
common.button.yes.label = Ja
common.button.no.label = Nej

common.confirmation = Bekr�ftelse
common.information = Information

common.message.error.invalidFileName            = Filnamnet kan inte inneh�lla tecknet:
common.message.error.canNotListFilesInDirectory = Kan inte lista filer i katalog:

common.missing.value = inget v�rde