help.title = Hjälp
help.text = Information:\n\n \
            This window will be used to configure the JavaPEG application.\n\n \
            It is possible to either import an configuration from an previous\n \
            installation or to specify which language to use in the application.\n\n \
            In section 1 (Configuration Mode) must a selection be done, either\n \
            should \"No Import\" set to selected, then must a language in the\n \
            section 2 (Configuration) be selected.\n\n \
            If \"Import\" is selected in section 1, then there are two possibilities,\n \
            either to select a configuration file from the list \"Found configurations\n \
            in user home directory\" (if the current user has done any previous\n \
            installations of JavaPEG that are possible to import), or to find\n \
            installations in another place by clicking the \"Import configuration from\n \
            other installation, select a directory in the directory selector that opens\n \
            and the select a configuration in the \"Found Configurations\" list.\n\n \
            When selections are done, then click the \"Continue\" button or the\n \
            \"Cancel\" button to abort the application configuration and start.

configuration.mode.title = 1: Konfigurations läge
configuration.mode.noimport = Ingen import
configuration.mode.import = Import

configuration.section.title = 2: Konfiguration
configuration.section.available.languages = Välj applikationsspråk:
configuration.section.available.configurations.in.user.home = Funna konfigurationer i användarens hemkatalog

configuration.section.other.import.location.title = Importera konfiguration från annan installation:
configuration.section.other.import.location.found.configurations = Funna konfigurationer