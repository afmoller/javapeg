category.categoriesModel.create.error = Kan inte ladda kategorier.\nJavaPEG kommer att avslutas\n\nSe loggfil f�r detaljer.
category.categoriesModel.store.error  = Kan inte spara kategorier.\nJavaPEG kommer att avslutas\n\nSe loggfil f�r detaljer.

category.categoriesModel.repositoryExists       = Bilddatabass�kv�g existerar.
category.categoriesModel.repositoryNotExists    = Bilddatabass�kv�g existerar inte.
category.categoriesModel.repositoryNotAvailable = Bilddatabass�kv�g inte tillg�nglig.

category.metadatavalue.selection.mode   = URVALSMETOD
category.metadatavalue.selection.values = V�RDEN

category.enterNameForNewCategory    = Please enter a name for the new category
category.enterNameForNewSubCategory = Please enter a name for the sub category

category.errormessage.categoryNameCanNotStartWithSpace = The category name can not start with a white space:
category.errormessage.categoryNameAlreadyExistsInScope = already exists as a category in the selected scope, please choose another name