# This is the Swedish language file for the category strings.

# The structure of the file is as follows:

# A line starting with "#" is interpreted as a comment.

# A valid non comment line may look like "file = Arkiv" where "file" is the variable, = the
# separator and "Arkiv" is the value of the variable, in this case the Swedish word for file.

# There might be whitespaces or tabs in between the variable and the "=". Any whitespace
# or other character after the value of the variable will be trimmed away.

# For more information regarding the rules for the syntax of this file please visit:
# http://java.sun.com/javase/6/docs/api/java/util/Properties.html

category.categoriesModel.create.error = Kan inte ladda kategorier.\nJavaPEG kommer att avslutas\n\nSe loggfil för detaljer.
category.categoriesModel.store.error  = Kan inte spara kategorier.\nJavaPEG kommer att avslutas\n\nSe loggfil för detaljer.

category.metadatavalue.selection.mode   = URVALSMETOD
category.metadatavalue.selection.values = VÄRDEN

category.enterNameForNewCategory    = Ange ett namn för den nya kategorin
category.enterNameForNewSubCategory = Ange ett namn för den nya underkategorin
category.enterNewNameForCategory    = Ange ett nytt namn för den kategorin:
category.rename                     = Byt namn på kategori

category.errormessage.categoryNameCanNotStartWithSpace = Kategorinamnet kan inte börja med ett mellanslag:
category.errormessage.categoryNameAlreadyExistsInScope = existerar redan som en kategori i vald kontext, välj ett annat namn

category.addToImageRepositoryHeader = Lägg till bild(er) till bilddatabas?
category.addToImageRepositoryQuestionPartOne = Lägg till bild(erna) i katalog:
category.addToImageRepositoryQuestionPartTwo = till bilddatabasen?

category.rememberMySelection = Kom ihåg mitt val (Kan ändras i Inställningarna)

category.mineCategoriesTab = Mina