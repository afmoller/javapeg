category.categoriesModel.create.error = Kan inte ladda kategorier.\nJavaPEG kommer att avslutas\n\nSe loggfil f�r detaljer.
category.categoriesModel.store.error