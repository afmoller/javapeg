category.categoriesModel.create.error = Kan inte ladda kategorier.\nJavaPEG kommer att avslutas\n\nSe loggfil f�r detaljer.
category.categoriesModel.store.error  = Kan inte spara kategorier.\nJavaPEG kommer att avslutas\n\nSe loggfil f�r detaljer.

category.categoriesModel.repositoryExists       = Bilddatabass�kv�g existerar.
category.categoriesModel.repositoryNotExists    = Bilddatabass�kv�g existerar inte.
category.categoriesModel.repositoryNotAvailable = Bilddatabass�kv�g inte tillg�nglig.