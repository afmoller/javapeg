category.categoriesModel.create.error = Kan inte ladda kategorier.\nJavaPEG kommer att avslutas\n\nSe loggfil f�r detaljer.
category.categoriesModel.store.error  = Kan inte spara kategorier.\nJavaPEG kommer att avslutas\n\nSe loggfil f�r detaljer.

category.categoriesModel.repositoryExists       = Bilddatabass�kv�g existerar.
category.categoriesModel.repositoryNotExists    = Bilddatabass�kv�g existerar inte.
category.categoriesModel.repositoryNotAvailable = Bilddatabass�kv�g inte tillg�nglig.

category.metadatavalue.selection.mode   = URVALSMETOD
category.metadatavalue.selection.values = V�RDEN

category.enterNameForNewCategory    = Ange ett namn f�r den nya kategorin
category.enterNameForNewSubCategory = Ange ett namn f�r den nya underkategorin
category.enterNewNameForCategory    = Ange ett nytt namn f�r den kategorin:
categrory.rename                    = Byt namn p� kategori

category.errormessage.categoryNameCanNotStartWithSpace = Kategorinamnet kan inte b�rja med ett mellanslag:
category.errormessage.categoryNameAlreadyExistsInScope = existerar redan som en kategori i vald kontext, v�lj ett annat namn

category.addToImageRepositoryHeader = L�gg till bild(er) till bilddatabas?
category.addToImageRepositoryQuestionPartOne = L�gg till bild(erna) i katalog:
category.addToImageRepositoryQuestionPartTwo = till bilddatabasen?