# This is the Swedish language file for the Image resizer part of JavaPEG.

# The structure of the file is as follows:

# A line starting with "#" is interpreted as a comment.

# A valid non comment line may look like "file = Arkiv" where "file" is the variable, = the
# separator and "Arkiv" is the value of the variable, in this case the Swedish word for file.

# There might be whitespaces or tabs in between the variable and the "=". Any whitespace
# or other character after the value of the variable will be trimmed away.

# For more information regarding the rules for the syntax of this file please visit:
# http://java.sun.com/javase/6/docs/api/java/util/Properties.html

imageresizer.gui.title = Bildstorleksändrare

imageresizer.processlog.title = PROCESSLOGG
imageresizer.processlog.image.processed = Bild: %s storleksändrad (%s) millisekunder)
imageresizer.processlog.image.resize.done = Storleksändringsprocessen tog: %s sekunder
imageresizer.processlog.image.resize.done.cancelled = Storleksändringsprocessen avbruten efter: %s sekunder

imageresizer.resize.input.width           = Bredd
imageresizer.resize.input.height          = Höjd
imageresizer.resize.input.keepaspectratio = Begränsande ram
imageresizer.resize.input.quality         = Kvalitet
imageresizer.resize.input.path            = Målkatalog

imageresizer.resize.input.button.resize = Storleksändra
imageresizer.resize.input.button.cancel = Avbryt

imageresizer.resize.process.destination.directory.created = Destinationskatalog skapad:
imageresizer.resize.process.couldNotCreateDirectory       = Kunde inte skapa katalog
imageresizer.resize.process.started                       = Storleksändringsprocess startad
imageresizer.resize.process.aborted                       = Storleksändringsprocess avbruten
imageresizer.resize.process.cancelled                     = Storleksändring avbruten
imageresizer.resize.process.done                          = Storleksändring färdig